-- THE REGISTERS IN VHDL
