---------------------------------------------------------------------
-- Control Unit
---------------------------------------------------------------------