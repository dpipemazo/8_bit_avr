---------------------------------------------------------------------
-- Memory Management Unit
---------------------------------------------------------------------