-- THE ALU
